module OBUF (
    input  I,
    output O
);
    assign O = I;
endmodule

