module VCC (
    output P
);
    assign P = 1'b1;
endmodule

