module IBUF (
    input  I,
    output O
);
    assign O = I;
endmodule

